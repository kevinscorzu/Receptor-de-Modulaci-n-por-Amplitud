module Adder (input logic [63:0] A, B,
				  output logic [63:0] C);
				
	assign C = A + B;
				
endmodule 