module Adder (input logic [31:0] A, B,
				  output logic [31:0] C);
				
	assign C = A + B;
				
endmodule 